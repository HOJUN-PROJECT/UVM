`include "fulladd10_en.v"
